`timescale 1ns / 1ps

module interface(

    );
endmodule
